module disp_ctrl 
# (
    parameter BIT_WIDTH = 20
)
(
    input logic [3:0] sel,
    output logic [0:BIT_WIDTH-1] bitmap [0:BIT_WIDTH-1]
);

always_comb begin : bitmap_block
    case (sel)
        4'h0: begin
            bitmap = '{
                20'b00000000111110000000,
                20'b00000001111111000000,
                20'b00000111111111110000,
                20'b00001111111111110000,
                20'b00001111111111111000,
                20'b00011111100011111000,
                20'b00011111000011111100,
                20'b00011111000011111100,
                20'b00011111000001111100,
                20'b00011111000001111100,
                20'b00011111000001111100,
                20'b00011111000001111100,
                20'b00011111000001111100,
                20'b00011111000011111100,
                20'b00011111000011111100,
                20'b00011111100111111000,
                20'b00001111111111111000,
                20'b00001111111111110000,
                20'b00000111111111110000,
                20'b00000001111111000000
            };
        end 
        4'h1: begin
            bitmap = '{
                20'b00000000000111110000,
                20'b00000000001111110000,
                20'b00000000011111110000,
                20'b00000000111111110000,
                20'b00000011111111110000,
                20'b00001111111111110000,
                20'b00001111111111110000,
                20'b00001111111111110000,
                20'b00001111001111110000,
                20'b00000000001111110000,
                20'b00000000001111110000,
                20'b00000000001111110000,
                20'b00000000001111110000,
                20'b00000000001111110000,
                20'b00000000001111110000,
                20'b00000000001111110000,
                20'b00000000001111110000,
                20'b00000000001111110000,
                20'b00000000001111110000,
                20'b00000000001111110000
            };
        end
        4'h2: begin
            bitmap = '{
                20'b00000001111111000000,
                20'b00000111111111110000,
                20'b00001111111111111000,
                20'b00001111111111111100,
                20'b00011111100011111100,
                20'b00011111100011111100,
                20'b00011111000011111100,
                20'b00000000000011111100,
                20'b00000000000111111000,
                20'b00000000001111111000,
                20'b00000000111111110000,
                20'b00000001111111100000,
                20'b00000011111110000000,
                20'b00000111111100000000,
                20'b00001111111000000000,
                20'b00001111111111111100,
                20'b00011111111111111100,
                20'b00011111111111111100,
                20'b00111111111111111100,
                20'b00111111111111111100
            };
        end 
        4'h3: begin
            bitmap = '{
                20'b00000000011100000000,
                20'b00000011111111100000,
                20'b00001111111111110000,
                20'b00001111111111111000,
                20'b00011111100111111000,
                20'b00011111000011111000,
                20'b00000000000111111000,
                20'b00000000001111110000,
                20'b00000000011111110000,
                20'b00000000011111110000,
                20'b00000000011111111000,
                20'b00000000000111111100,
                20'b00000000000011111100,
                20'b00000000000011111100,
                20'b00011111000011111100,
                20'b00011111100011111100,
                20'b00011111111111111000,
                20'b00001111111111111000,
                20'b00000111111111100000,
                20'b00000000111110000000
            };
        end 
        4'h4: begin
            bitmap = '{
                20'b00000000000001110000,
                20'b00000000000111110000,
                20'b00000000001111110000,
                20'b00000000011111110000,
                20'b00000000111111110000,
                20'b00000001111111110000,
                20'b00000001111111110000,
                20'b00000011111111110000,
                20'b00000111110111110000,
                20'b00001111100111110000,
                20'b00011111000111110000,
                20'b00111111000111110000,
                20'b00111111111111111100,
                20'b00111111111111111110,
                20'b00111111111111111110,
                20'b00111111111111111110,
                20'b00000000000111111000,
                20'b00000000000111110000,
                20'b00000000000111110000,
                20'b00000000000111110000
            };
        end 
        4'h5: begin
            bitmap = '{
                20'b00000111111111111000,
                20'b00000111111111111000,
                20'b00001111111111111000,
                20'b00001111111111111000,
                20'b00001111111111111000,
                20'b00001111100000000000,
                20'b00001111100000000000,
                20'b00001111111111100000,
                20'b00001111111111110000,
                20'b00011111111111111000,
                20'b00011111111111111100,
                20'b00000001000011111100,
                20'b00000000000011111100,
                20'b00000000000001111100,
                20'b00011111000001111100,
                20'b00011111100011111100,
                20'b00011111111111111000,
                20'b00001111111111111000,
                20'b00000111111111110000,
                20'b00000001111111000000
            };
        end 
        4'h6: begin
            bitmap = '{
                20'b00000000111110000000,
                20'b00000001111111000000,
                20'b00000111111111110000,
                20'b00001111111111111000,
                20'b00001111111111111000,
                20'b00011111100011111000,
                20'b00011111000000000000,
                20'b00011111000111000000,
                20'b00011111111111110000,
                20'b00111111111111111000,
                20'b00111111111111111000,
                20'b00111111100011111100,
                20'b00011111000011111100,
                20'b00011111000001111100,
                20'b00011111000001111100,
                20'b00011111100011111100,
                20'b00001111111111111000,
                20'b00001111111111111000,
                20'b00000111111111110000,
                20'b00000001111111000000
            };
        end 
        4'h7: begin
            bitmap = '{
                20'b00111111111111111100,
                20'b00111111111111111100,
                20'b00111111111111111100,
                20'b00111111111111111100,
                20'b00011111111111111000,
                20'b00000000000111110000,
                20'b00000000001111100000,
                20'b00000000011111100000,
                20'b00000000011111000000,
                20'b00000000111111000000,
                20'b00000000111110000000,
                20'b00000001111110000000,
                20'b00000001111100000000,
                20'b00000001111100000000,
                20'b00000011111100000000,
                20'b00000011111000000000,
                20'b00000011111000000000,
                20'b00000011111000000000,
                20'b00000011111000000000,
                20'b00000011111000000000
            };
        end 
        4'h8: begin
            bitmap = '{
                20'b00000001111110000000,
                20'b00000111111111100000,
                20'b00001111111111110000,
                20'b00011111111111111000,
                20'b00011111100011111000,
                20'b00011111000011111000,
                20'b00011111100111111000,
                20'b00001111111111110000,
                20'b00000111111111110000,
                20'b00001111111111110000,
                20'b00011111111111111000,
                20'b00011111100111111000,
                20'b00011111000011111100,
                20'b00011111000011111100,
                20'b00011111000011111100,
                20'b00011111100111111000,
                20'b00011111111111111000,
                20'b00001111111111110000,
                20'b00000111111111100000,
                20'b00000000111110000000
            };
        end 
        4'h9: begin
            bitmap = '{
                20'b00000000111000000000,
                20'b00000111111111000000,
                20'b00001111111111100000,
                20'b00011111111111110000,
                20'b00011111100111111000,
                20'b00011111000011111000,
                20'b00111111000011111000,
                20'b00111111000011111100,
                20'b00011111000011111100,
                20'b00011111100111111100,
                20'b00011111111111111100,
                20'b00001111111111111100,
                20'b00000111111011111100,
                20'b00000000000011111000,
                20'b00000011000011111000,
                20'b00011111100111111000,
                20'b00011111111111110000,
                20'b00001111111111110000,
                20'b00000111111111000000,
                20'b00000001111100000000
            };
        end 
        default: begin
                        bitmap = '{
                20'b00000001111001111000,
                20'b00000001111001111000,
                20'b00000001110001111000,
                20'b00000011110001111000,
                20'b00000011110011110000,
                20'b00011111111111111100,
                20'b00111111111111111100,
                20'b00111111111111111100,
                20'b00011111111111111100,
                20'b00000111100111100000,
                20'b00000111100111100000,
                20'b00000111100111100000,
                20'b00011111111111111100,
                20'b00111111111111111100,
                20'b00111111111111111100,
                20'b00011111111111100000,
                20'b00001111001111000000,
                20'b00001111001111000000,
                20'b00011110001111000000,
                20'b00011110001111000000
            };
        end
    endcase
end
endmodule